library verilog;
use verilog.vl_types.all;
entity ALU_4_vlg_vec_tst is
end ALU_4_vlg_vec_tst;
