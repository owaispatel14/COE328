library verilog;
use verilog.vl_types.all;
entity ModifiedControlUnit_vlg_vec_tst is
end ModifiedControlUnit_vlg_vec_tst;
